`timescale 1ns / 1ps

module systolicarray_2_tb(

    );

parameter size=8;
parameter decimal=4;

reg clk,rst;
reg[4*size-1:0] mi0;
reg[4*size-1:0] mi1;
wire[4*size-1:0] mor;

systolicarray_2 s2(clk,rst,mi0,mi1,mor);

initial begin
clk=0;
rst=0;
//  |0.5 1 |   |1 2|
//  |1  0.5| x |3 4|  
mi0=8|(16<<8)|(16<<16)|(8<<24);     //  mi0 = [8][16][16][8] = [0.5][1][1][0.5].
mi1=16|(32<<8)|(48<<16)|(64<<24);   //  mi1 = [16][31][48][64] = [1][2][3][4].

#4 rst=1;

end

always #1 begin
    clk<=~clk;
end

endmodule
